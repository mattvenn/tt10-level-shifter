magic
tech sky130A
magscale 1 2
timestamp 1740491262
<< pwell >>
rect -256 -221 256 221
<< nmos >>
rect -60 -11 60 73
<< ndiff >>
rect -118 61 -60 73
rect -118 1 -106 61
rect -72 1 -60 61
rect -118 -11 -60 1
rect 60 61 118 73
rect 60 1 72 61
rect 106 1 118 61
rect 60 -11 118 1
<< ndiffc >>
rect -106 1 -72 61
rect 72 1 106 61
<< psubdiff >>
rect -220 151 -124 185
rect 124 151 220 185
rect -220 89 -186 151
rect 186 89 220 151
rect -220 -151 -186 -89
rect 186 -151 220 -89
rect -220 -185 -124 -151
rect 124 -185 220 -151
<< psubdiffcont >>
rect -124 151 124 185
rect -220 -89 -186 89
rect 186 -89 220 89
rect -124 -185 124 -151
<< poly >>
rect -60 73 60 99
rect -60 -49 60 -11
rect -60 -83 -44 -49
rect 44 -83 60 -49
rect -60 -99 60 -83
<< polycont >>
rect -44 -83 44 -49
<< locali >>
rect -220 151 -124 185
rect 124 151 220 185
rect -220 89 -186 151
rect 186 89 220 151
rect -106 61 -72 77
rect -106 -15 -72 1
rect 72 61 106 77
rect 72 -15 106 1
rect -60 -83 -44 -49
rect 44 -83 60 -49
rect -220 -151 -186 -89
rect 186 -151 220 -89
rect -220 -185 -124 -151
rect 124 -185 220 -151
<< viali >>
rect -106 1 -72 61
rect 72 1 106 61
rect -44 -83 44 -49
<< metal1 >>
rect -112 61 -66 73
rect -112 1 -106 61
rect -72 1 -66 61
rect -112 -11 -66 1
rect 66 61 112 73
rect 66 1 72 61
rect 106 1 112 61
rect 66 -11 112 1
rect -56 -49 56 -43
rect -56 -83 -44 -49
rect 44 -83 56 -49
rect -56 -89 56 -83
<< properties >>
string FIXED_BBOX -203 -168 203 168
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.6 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
