magic
tech sky130A
magscale 1 2
timestamp 1740491448
<< error_p >>
rect -29 -179 29 -173
rect -29 -213 -17 -179
rect -29 -219 29 -213
<< nwell >>
rect -226 -352 226 352
<< pmoshvt >>
rect -30 -132 30 204
<< pdiff >>
rect -88 192 -30 204
rect -88 -120 -76 192
rect -42 -120 -30 192
rect -88 -132 -30 -120
rect 30 192 88 204
rect 30 -120 42 192
rect 76 -120 88 192
rect 30 -132 88 -120
<< pdiffc >>
rect -76 -120 -42 192
rect 42 -120 76 192
<< nsubdiff >>
rect -190 282 -94 316
rect 94 282 190 316
rect -190 219 -156 282
rect 156 219 190 282
rect -190 -282 -156 -219
rect 156 -282 190 -219
rect -190 -316 -94 -282
rect 94 -316 190 -282
<< nsubdiffcont >>
rect -94 282 94 316
rect -190 -219 -156 219
rect 156 -219 190 219
rect -94 -316 94 -282
<< poly >>
rect -30 204 30 230
rect -30 -163 30 -132
rect -33 -179 33 -163
rect -33 -213 -17 -179
rect 17 -213 33 -179
rect -33 -229 33 -213
<< polycont >>
rect -17 -213 17 -179
<< locali >>
rect -190 282 -94 316
rect 94 282 190 316
rect -190 219 -156 282
rect 156 219 190 282
rect -76 192 -42 208
rect -76 -136 -42 -120
rect 42 192 76 208
rect 42 -136 76 -120
rect -33 -213 -17 -179
rect 17 -213 33 -179
rect -190 -282 -156 -219
rect 156 -282 190 -219
rect -190 -316 -94 -282
rect 94 -316 190 -282
<< viali >>
rect -76 -120 -42 192
rect 42 -120 76 192
rect -17 -213 17 -179
<< metal1 >>
rect -82 192 -36 204
rect -82 -120 -76 192
rect -42 -120 -36 192
rect -82 -132 -36 -120
rect 36 192 82 204
rect 36 -120 42 192
rect 76 -120 82 192
rect 36 -132 82 -120
rect -29 -179 29 -173
rect -29 -213 -17 -179
rect 17 -213 29 -179
rect -29 -219 29 -213
<< properties >>
string FIXED_BBOX -173 -299 173 299
string gencell sky130_fd_pr__pfet_01v8_hvt
string library sky130
string parameters w 1.68 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
