magic
tech sky130A
magscale 1 2
timestamp 1740492959
<< pwell >>
rect 5620 -300 5820 -100
rect 5760 -1240 6200 -1180
rect 5200 -1360 5380 -1340
rect 5200 -1420 5400 -1360
rect 4520 -1540 4580 -1460
rect 5340 -1540 5400 -1420
<< viali >>
rect 4800 -540 4980 -500
rect 5220 -540 5400 -500
rect 5640 -540 5820 -500
rect 6080 -680 6260 -640
rect 3660 -780 3820 -740
rect 4380 -800 4540 -760
rect 3660 -1680 3820 -1640
rect 4380 -1660 4560 -1620
rect 5240 -1660 5420 -1620
rect 5660 -1660 5840 -1620
rect 6100 -1660 6280 -1620
<< metal1 >>
rect 3520 -740 3940 -100
rect 3520 -780 3660 -740
rect 3820 -780 3940 -740
rect 3520 -800 3940 -780
rect 4220 -360 5060 -100
rect 5620 -200 5820 -100
rect 5620 -220 5960 -200
rect 5620 -300 5860 -220
rect 5940 -300 5960 -220
rect 4220 -500 6380 -360
rect 4220 -540 4800 -500
rect 4980 -540 5220 -500
rect 5400 -540 5640 -500
rect 5820 -540 6380 -500
rect 4220 -560 6380 -540
rect 4220 -760 4660 -560
rect 4220 -800 4380 -760
rect 4540 -800 4660 -760
rect 3620 -960 3700 -800
rect 4220 -820 4660 -800
rect 3760 -1000 3820 -880
rect 4340 -960 4400 -820
rect 4480 -960 4600 -880
rect 4780 -960 4840 -560
rect 4920 -780 5000 -620
rect 5680 -660 5700 -600
rect 5760 -660 5780 -600
rect 5960 -640 6380 -560
rect 5960 -680 6080 -640
rect 6260 -680 6380 -640
rect 5960 -720 6380 -680
rect 4920 -800 5040 -780
rect 4920 -860 4960 -800
rect 5020 -860 5040 -800
rect 4920 -880 5040 -860
rect 4920 -960 5000 -880
rect 5180 -940 5280 -720
rect 5340 -800 5700 -720
rect 5340 -860 5500 -800
rect 5560 -860 5700 -800
rect 5340 -940 5700 -860
rect 5180 -960 5260 -940
rect 4560 -1000 4600 -960
rect 3700 -1180 3820 -1000
rect 4040 -1180 4160 -1160
rect 3700 -1260 4060 -1180
rect 4140 -1260 4160 -1180
rect 3700 -1380 3820 -1260
rect 4040 -1280 4160 -1260
rect 4400 -1180 4520 -1000
rect 4560 -1060 4940 -1000
rect 4560 -1180 4600 -1060
rect 4400 -1260 4600 -1180
rect 3700 -1440 3880 -1380
rect 4400 -1420 4520 -1260
rect 3620 -1600 3700 -1480
rect 3800 -1560 3880 -1440
rect 4320 -1600 4380 -1440
rect 4560 -1460 4600 -1260
rect 5180 -1140 5240 -960
rect 5280 -1020 5380 -1000
rect 5280 -1080 5300 -1020
rect 5360 -1080 5380 -1020
rect 5280 -1100 5380 -1080
rect 5180 -1340 5260 -1140
rect 5760 -1180 5820 -800
rect 6080 -940 6140 -720
rect 6180 -920 6500 -780
rect 6100 -1180 6200 -980
rect 5760 -1240 6200 -1180
rect 5180 -1360 5380 -1340
rect 5180 -1420 5800 -1360
rect 4520 -1540 4600 -1460
rect 4840 -1600 5040 -1480
rect 5200 -1600 5260 -1460
rect 5340 -1540 5400 -1420
rect 5860 -1460 5940 -1240
rect 6100 -1420 6200 -1240
rect 6400 -1020 6500 -920
rect 6400 -1220 6640 -1020
rect 6400 -1460 6500 -1220
rect 5640 -1600 5700 -1460
rect 5780 -1520 5940 -1460
rect 6080 -1600 6140 -1460
rect 6200 -1520 6500 -1460
rect 3500 -1620 6380 -1600
rect 3500 -1640 4380 -1620
rect 3500 -1680 3660 -1640
rect 3820 -1660 4380 -1640
rect 4560 -1660 5240 -1620
rect 5420 -1660 5660 -1620
rect 5840 -1660 6100 -1620
rect 6280 -1660 6380 -1620
rect 3820 -1680 6380 -1660
rect 3500 -1820 6380 -1680
<< via1 >>
rect 5860 -300 5940 -220
rect 5700 -660 5760 -600
rect 4960 -860 5020 -800
rect 5500 -860 5560 -800
rect 4060 -1260 4140 -1180
rect 5300 -1080 5360 -1020
<< metal2 >>
rect 5840 -220 5960 -200
rect 5840 -300 5860 -220
rect 5940 -300 5960 -220
rect 5840 -600 5960 -300
rect 5680 -660 5700 -600
rect 5760 -660 5960 -600
rect 5680 -680 5960 -660
rect 4940 -800 5580 -780
rect 4940 -860 4960 -800
rect 5020 -860 5500 -800
rect 5560 -860 5580 -800
rect 4940 -880 5580 -860
rect 5280 -1020 5380 -1000
rect 5280 -1080 5300 -1020
rect 5360 -1080 5380 -1020
rect 5280 -1100 5380 -1080
rect 4040 -1180 4160 -1160
rect 5280 -1180 5360 -1100
rect 4040 -1260 4060 -1180
rect 4140 -1260 5360 -1180
rect 4040 -1280 4160 -1260
use sky130_fd_pr__nfet_01v8_48YY59  sky130_fd_pr__nfet_01v8_48YY59_0
timestamp 1740491262
transform 1 0 4456 0 -1 -1459
box -256 -221 256 221
use sky130_fd_pr__nfet_01v8_L6RDF9  sky130_fd_pr__nfet_01v8_L6RDF9_0
timestamp 1740491448
transform 1 0 5746 0 1 -1459
box -226 -221 226 221
use sky130_fd_pr__pfet_01v8_hvt_MY4TMJ  sky130_fd_pr__pfet_01v8_hvt_MY4TMJ_0
timestamp 1740491919
transform 1 0 5731 0 1 -828
box -211 -352 211 352
use sky130_fd_pr__pfet_01v8_hvt_GCT3R5  XM1
timestamp 1740491448
transform 1 0 4886 0 1 -828
box -226 -352 226 352
use sky130_fd_pr__pfet_01v8_hvt_6W9GZD  XM2
timestamp 1740491448
transform 1 0 4446 0 1 -954
box -226 -226 226 226
use sky130_fd_pr__pfet_01v8_hvt_M479BK  XM4
timestamp 1740491262
transform 1 0 3731 0 -1 -954
box -211 -226 211 226
use sky130_fd_pr__pfet_01v8_hvt_LY4TMQ  XM5
timestamp 1740491448
transform 1 0 5311 0 1 -828
box -211 -352 211 352
use sky130_fd_pr__nfet_01v8_L6RDF9  XM7
timestamp 1740491448
transform 1 0 5306 0 1 -1459
box -226 -221 226 221
use sky130_fd_pr__nfet_01v8_L78EGD  XM9
timestamp 1740491448
transform 1 0 6171 0 1 -1459
box -211 -221 211 221
use sky130_fd_pr__pfet_01v8_hvt_2MG8BZ  XM10
timestamp 1740491448
transform 1 0 6151 0 1 -892
box -211 -268 211 268
use sky130_fd_pr__nfet_01v8_48YY59  XM11
timestamp 1740491262
transform 1 0 3757 0 -1 -1478
box -256 -221 256 221
<< labels >>
flabel metal1 4800 -300 5000 -100 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 4840 -1680 5040 -1480 0 FreeSans 256 0 0 0 GND
port 0 nsew
flabel metal1 3640 -300 3840 -100 0 FreeSans 256 0 0 0 VDD_L
port 2 nsew
flabel metal1 3740 -1260 4140 -1180 0 FreeSans 400 0 0 0 src_n
flabel metal1 6440 -1220 6640 -1020 0 FreeSans 256 0 0 0 OUT
port 4 nsew
flabel metal1 6100 -1420 6200 -980 0 FreeSans 400 0 0 0 out_n
flabel metal1 5620 -300 5820 -100 0 FreeSans 256 0 0 0 IN
port 3 nsew
flabel space 5200 -1420 5260 -720 0 FreeSans 400 0 0 0 out_p
flabel metal1 4560 -1060 4940 -1000 0 FreeSans 400 0 0 0 net2
flabel metal2 5020 -880 5500 -780 0 FreeSans 400 0 0 0 net1
<< end >>
