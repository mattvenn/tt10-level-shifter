magic
tech sky130A
magscale 1 2
timestamp 1740499851
<< viali >>
rect 18300 42730 18340 42770
rect 18410 42730 18450 42770
<< metal1 >>
rect 17874 43020 17880 43140
rect 18000 43020 18560 43140
rect 18280 42770 18360 42790
rect 17960 42760 18020 42766
rect 18280 42760 18300 42770
rect 18020 42730 18300 42760
rect 18340 42730 18360 42770
rect 18020 42700 18360 42730
rect 18390 42770 18500 42790
rect 18390 42730 18410 42770
rect 18450 42760 18500 42770
rect 18450 42730 20340 42760
rect 18390 42720 20340 42730
rect 18390 42710 18500 42720
rect 17960 42694 18020 42700
rect 16480 42420 18560 42540
rect 16480 41040 16600 42420
rect 19020 42080 19220 42086
rect 18276 41742 18282 41898
rect 18438 41742 18444 41898
rect 19220 41880 19460 42080
rect 19020 41874 19220 41880
rect 18282 41442 18438 41742
rect 19260 41460 19460 41880
rect 20300 41580 20340 42720
rect 16480 40914 16600 40920
rect 21220 40580 21390 40640
rect 21450 40580 21456 40640
rect 17920 40120 18260 40160
rect 17920 39940 17940 40120
rect 18100 39960 18324 40120
rect 18100 39940 18260 39960
rect 17920 39900 18260 39940
<< via1 >>
rect 17880 43020 18000 43140
rect 17960 42700 18020 42760
rect 18282 41742 18438 41898
rect 19020 41880 19220 42080
rect 16480 40920 16600 41040
rect 21390 40580 21450 40640
rect 17940 39940 18100 40120
<< metal2 >>
rect 17880 43140 18000 43146
rect 17511 43020 17520 43140
rect 17640 43020 17880 43140
rect 17880 43014 18000 43020
rect 17872 42760 17928 42767
rect 17870 42758 17960 42760
rect 17870 42702 17872 42758
rect 17928 42702 17960 42758
rect 17870 42700 17960 42702
rect 18020 42700 18026 42760
rect 17872 42693 17928 42700
rect 17207 42598 17353 42602
rect 17202 42593 17358 42598
rect 17202 42447 17207 42593
rect 17353 42447 17358 42593
rect 17202 42318 17358 42447
rect 17202 42162 18438 42318
rect 18282 41898 18438 42162
rect 18845 42080 19035 42084
rect 18840 42075 19020 42080
rect 18840 41885 18845 42075
rect 18840 41880 19020 41885
rect 19220 41880 19226 42080
rect 18845 41876 19035 41880
rect 18282 41736 18438 41742
rect 16474 40920 16480 41040
rect 16600 40920 16606 41040
rect 16480 40860 16600 40920
rect 16480 40731 16600 40740
rect 21390 40640 21450 40646
rect 21450 40580 21680 40640
rect 21390 40574 21450 40580
rect 21620 40208 21680 40580
rect 17500 40140 18140 40160
rect 21613 40152 21622 40208
rect 21678 40152 21687 40208
rect 21620 40150 21680 40152
rect 17500 39920 17520 40140
rect 17740 40120 18140 40140
rect 17740 39940 17940 40120
rect 18100 39940 18140 40120
rect 17740 39920 18140 39940
rect 17500 39900 18140 39920
<< via2 >>
rect 17520 43020 17640 43140
rect 17872 42702 17928 42758
rect 17207 42447 17353 42593
rect 18845 41885 19020 42075
rect 19020 41885 19035 42075
rect 16480 40740 16600 40860
rect 21622 40152 21678 40208
rect 17520 39920 17740 40140
<< metal3 >>
rect 1320 43180 17450 43200
rect 1320 42930 1430 43180
rect 1770 43140 17450 43180
rect 17515 43140 17645 43145
rect 1770 43020 17520 43140
rect 17640 43020 17645 43140
rect 1770 42930 17450 43020
rect 17515 43015 17645 43020
rect 1320 42900 17450 42930
rect 17202 42593 17358 42900
rect 17728 42762 17792 42768
rect 17867 42760 17933 42763
rect 17792 42758 17933 42760
rect 17792 42702 17872 42758
rect 17928 42702 17933 42758
rect 17792 42700 17933 42702
rect 17728 42692 17792 42698
rect 17867 42697 17933 42700
rect 17202 42447 17207 42593
rect 17353 42447 17358 42593
rect 17202 42442 17358 42447
rect 17640 42075 19040 42080
rect 17640 41885 18845 42075
rect 19035 41885 19040 42075
rect 17640 41880 19040 41885
rect 17640 41830 17960 41880
rect 200 41790 17960 41830
rect 200 41420 240 41790
rect 570 41420 17960 41790
rect 200 41390 17960 41420
rect 16475 40860 16605 40865
rect 16475 40740 16480 40860
rect 16600 40740 16605 40860
rect 16475 40735 16605 40740
rect 16480 40170 16600 40735
rect 21617 40208 21683 40213
rect 770 40140 17770 40170
rect 21617 40152 21622 40208
rect 21678 40152 21683 40208
rect 21617 40147 21683 40152
rect 770 39910 840 40140
rect 1180 39920 17520 40140
rect 17740 39920 17770 40140
rect 1180 39910 17770 39920
rect 770 39890 17770 39910
rect 21620 39542 21680 40147
rect 21612 39478 21618 39542
rect 21682 39478 21688 39542
<< via3 >>
rect 1430 42930 1770 43180
rect 17728 42698 17792 42762
rect 240 41420 570 41790
rect 840 39910 1180 40140
rect 21618 39478 21682 39542
<< metal4 >>
rect 3006 44952 3066 45152
rect 3558 44952 3618 45152
rect 4110 44952 4170 45152
rect 4662 44952 4722 45152
rect 5214 44952 5274 45152
rect 5766 44952 5826 45152
rect 6318 44952 6378 45152
rect 6870 44952 6930 45152
rect 7422 44952 7482 45152
rect 7974 44952 8034 45152
rect 8526 44952 8586 45152
rect 9078 44952 9138 45152
rect 9630 44952 9690 45152
rect 10182 44952 10242 45152
rect 10734 44952 10794 45152
rect 11286 44952 11346 45152
rect 11838 44952 11898 45152
rect 12390 44952 12450 45152
rect 12942 44952 13002 45152
rect 13494 44952 13554 45152
rect 14046 44952 14106 45152
rect 14598 44952 14658 45152
rect 15150 44952 15210 45152
rect 200 41790 600 44152
rect 200 41420 240 41790
rect 570 41420 600 41790
rect 200 1000 600 41420
rect 800 40140 1200 44152
rect 800 39910 840 40140
rect 1180 39910 1200 40140
rect 800 1000 1200 39910
rect 1400 43180 1800 44152
rect 1400 42930 1430 43180
rect 1770 42930 1800 43180
rect 1400 1000 1800 42930
rect 15702 39540 15762 45152
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 44952 20730 45152
rect 21222 44952 21282 45152
rect 21774 44952 21834 45152
rect 22326 44952 22386 45152
rect 22878 44952 22938 45152
rect 23430 44952 23490 45152
rect 23982 44952 24042 45152
rect 24534 43590 24594 45152
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 17730 43530 24594 43590
rect 17730 42763 17790 43530
rect 17727 42762 17793 42763
rect 17727 42698 17728 42762
rect 17792 42698 17793 42762
rect 17727 42697 17793 42698
rect 21617 39542 21683 39543
rect 21617 39540 21618 39542
rect 15702 39480 21618 39540
rect 21617 39478 21618 39480
rect 21682 39478 21683 39542
rect 21617 39477 21683 39478
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 27234 0 27414 200
use level_shifter2  level_shifter2_0
timestamp 1740494155
transform 1 0 14664 0 1 41766
box 3500 -1820 6640 -100
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0
timestamp 1704896540
transform 1 0 18278 0 1 42508
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1704896540
transform 1 0 18188 0 1 42508
box -38 -48 130 592
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 1400 1000 1800 44152 1 FreeSans 1600 0 0 0 VAPWR
port 53 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
