magic
tech sky130A
magscale 1 2
timestamp 1740491448
<< error_p >>
rect -29 83 29 89
rect -29 49 -17 83
rect -29 43 29 49
<< pwell >>
rect -226 -221 226 221
<< nmos >>
rect -30 -73 30 11
<< ndiff >>
rect -88 -1 -30 11
rect -88 -61 -76 -1
rect -42 -61 -30 -1
rect -88 -73 -30 -61
rect 30 -1 88 11
rect 30 -61 42 -1
rect 76 -61 88 -1
rect 30 -73 88 -61
<< ndiffc >>
rect -76 -61 -42 -1
rect 42 -61 76 -1
<< psubdiff >>
rect -190 151 -94 185
rect 94 151 190 185
rect -190 89 -156 151
rect 156 89 190 151
rect -190 -151 -156 -89
rect 156 -151 190 -89
rect -190 -185 -94 -151
rect 94 -185 190 -151
<< psubdiffcont >>
rect -94 151 94 185
rect -190 -89 -156 89
rect 156 -89 190 89
rect -94 -185 94 -151
<< poly >>
rect -33 83 33 99
rect -33 49 -17 83
rect 17 49 33 83
rect -33 33 33 49
rect -30 11 30 33
rect -30 -99 30 -73
<< polycont >>
rect -17 49 17 83
<< locali >>
rect -190 151 -94 185
rect 94 151 190 185
rect -190 89 -156 151
rect 156 89 190 151
rect -33 49 -17 83
rect 17 49 33 83
rect -76 -1 -42 15
rect -76 -77 -42 -61
rect 42 -1 76 15
rect 42 -77 76 -61
rect -190 -151 -156 -89
rect 156 -151 190 -89
rect -190 -185 -94 -151
rect 94 -185 190 -151
<< viali >>
rect -17 49 17 83
rect -76 -61 -42 -1
rect 42 -61 76 -1
<< metal1 >>
rect -29 83 29 89
rect -29 49 -17 83
rect 17 49 29 83
rect -29 43 29 49
rect -82 -1 -36 11
rect -82 -61 -76 -1
rect -42 -61 -36 -1
rect -82 -73 -36 -61
rect 36 -1 82 11
rect 36 -61 42 -1
rect 76 -61 82 -1
rect 36 -73 82 -61
<< properties >>
string FIXED_BBOX -173 -168 173 168
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
