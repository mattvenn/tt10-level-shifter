magic
tech sky130A
magscale 1 2
timestamp 1740491448
<< error_p >>
rect -29 -179 29 -173
rect -29 -213 -17 -179
rect -29 -219 29 -213
<< nwell >>
rect -211 -352 211 352
<< pmoshvt >>
rect -15 -132 15 204
<< pdiff >>
rect -73 192 -15 204
rect -73 -120 -61 192
rect -27 -120 -15 192
rect -73 -132 -15 -120
rect 15 192 73 204
rect 15 -120 27 192
rect 61 -120 73 192
rect 15 -132 73 -120
<< pdiffc >>
rect -61 -120 -27 192
rect 27 -120 61 192
<< nsubdiff >>
rect -175 282 -79 316
rect 79 282 175 316
rect -175 219 -141 282
rect 141 219 175 282
rect -175 -282 -141 -219
rect 141 -282 175 -219
rect -175 -316 -79 -282
rect 79 -316 175 -282
<< nsubdiffcont >>
rect -79 282 79 316
rect -175 -219 -141 219
rect 141 -219 175 219
rect -79 -316 79 -282
<< poly >>
rect -15 204 15 230
rect -15 -163 15 -132
rect -33 -179 33 -163
rect -33 -213 -17 -179
rect 17 -213 33 -179
rect -33 -229 33 -213
<< polycont >>
rect -17 -213 17 -179
<< locali >>
rect -175 282 -79 316
rect 79 282 175 316
rect -175 219 -141 282
rect 141 219 175 282
rect -61 192 -27 208
rect -61 -136 -27 -120
rect 27 192 61 208
rect 27 -136 61 -120
rect -33 -213 -17 -179
rect 17 -213 33 -179
rect -175 -282 -141 -219
rect 141 -282 175 -219
rect -175 -316 -79 -282
rect 79 -316 175 -282
<< viali >>
rect -61 -120 -27 192
rect 27 -120 61 192
rect -17 -213 17 -179
<< metal1 >>
rect -67 192 -21 204
rect -67 -120 -61 192
rect -27 -120 -21 192
rect -67 -132 -21 -120
rect 21 192 67 204
rect 21 -120 27 192
rect 61 -120 67 192
rect 21 -132 67 -120
rect -29 -179 29 -173
rect -29 -213 -17 -179
rect 17 -213 29 -179
rect -29 -219 29 -213
<< properties >>
string FIXED_BBOX -158 -299 158 299
string gencell sky130_fd_pr__pfet_01v8_hvt
string library sky130
string parameters w 1.68 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
